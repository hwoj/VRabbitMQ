module vrabbitmq

fn main() {
	println('Hello World!')
}
